

module top(input clk)

endmodule
